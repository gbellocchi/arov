

/* =====================================================================
 * Project:      Accelerator-rich overlay
 * Title:        post_synth_tb_exilzcu102.sv
 * Description:  Post-synthesis testbench to launch related simulations
 *               for verification, power, etc.
 *
 * $Date:        26.7.2022
 * ===================================================================== */

`timescale 1 ps / 1 ps

module arov_tb();

  hero_exilzcu102 hero_exilzcu102_i();

endmodule